LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY SHIFT_OUT IS
	GENERIC (BIT_WIDTH : INTEGER := 8);
	PORT (CLK : IN STD_LOGIC;
			RST : IN STD_LOGIC;
			EN : IN STD_LOGIC;
			REG_IN : IN STD_LOGIC_VECTOR(BIT_WIDTH-1 DOWNTO 0);
			BIT_OUT : OUT STD_LOGIC);
END SHIFT_OUT;

ARCHITECTURE SHIFT_LOGIC OF SHIFT_OUT IS
	SIGNAL SHIFT_REGISTER : STD_LOGIC_VECTOR(BIT_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
BEGIN
	PROCESS(CLK, RST)
	BEGIN
		IF RST = '1' THEN
			SHIFT_REGISTER <= (OTHERS => '0');
		ELSIF CLK'EVENT AND CLK = '0' THEN
			IF EN = '0' THEN
				SHIFT_REGISTER <= SHIFT_REGISTER(BIT_WIDTH-2 DOWNTO 0) & '0';
			ELSE
				SHIFT_REGISTER(BIT_WIDTH-1 DOWNTO 0) <= REG_IN(BIT_WIDTH-1 DOWNTO 0);
			END IF;
		END IF;
	END PROCESS;
	BIT_OUT <= SHIFT_REGISTER(SHIFT_REGISTER'HIGH);
END SHIFT_LOGIC;
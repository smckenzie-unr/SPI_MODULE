LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY COUNTER IS
	GENERIC(BIT_WIDTH : INTEGER := 8);
	PORT(CLK : IN STD_LOGIC;
		  RST : IN STD_LOGIC;
		  EN : IN STD_LOGIC;
		  BITS_OUT : OUT STD_LOGIC_VECTOR(BIT_WIDTH-1 DOWNTO 0));
END COUNTER;

ARCHITECTURE LOGIC OF COUNTER IS
	SIGNAL COUNTER_REG : STD_LOGIC_VECTOR(BIT_WIDTH-1 DOWNTO 0);
BEGIN
	PROCESS(CLK, RST)
	BEGIN
		IF RST = '1' THEN
			COUNTER_REG <= (OTHERS => '0');
		ELSIF CLK'EVENT AND CLK = '1' THEN
			IF EN = '1' THEN
				COUNTER_REG <= COUNTER_REG + 1;
			END IF;
		END IF;
	END PROCESS;
	BITS_OUT(BIT_WIDTH-1 DOWNTO 0) <= COUNTER_REG(BIT_WIDTH-1 DOWNTO 0);
END LOGIC;
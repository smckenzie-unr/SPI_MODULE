LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY SPI_MODULE IS
	GENERIC(WORD_SIZE : INTEGER := 8);
	PORT(CLOCK : IN STD_LOGIC;
		  START_TRANSACTION : IN STD_LOGIC;
		  RESET_RX : IN STD_LOGIC;
		  REG_TX : IN STD_LOGIC_VECTOR(WORD_SIZE-1 DOWNTO 0);
		  MISO : IN STD_LOGIC;
		  REG_RX : OUT STD_LOGIC_VECTOR(WORD_SIZE-1 DOWNTO 0);
		  CHIP_SELECT : OUT STD_LOGIC;
		  MOSI : OUT STD_LOGIC);
END SPI_MODULE;

ARCHITECTURE BEHAVIOR OF SPI_MODULE IS
	COMPONENT SHIFT_IN IS
		GENERIC(BIT_WIDTH : INTEGER := WORD_SIZE);
		PORT(CLK : IN STD_LOGIC;
			  RST : IN STD_LOGIC;
			  EN : IN STD_LOGIC;
			  BIT_IN : IN STD_LOGIC;
			  REG_OUT : OUT STD_LOGIC_VECTOR(BIT_WIDTH-1 DOWNTO 0));
	END COMPONENT;
	COMPONENT SHIFT_OUT IS
		GENERIC(BIT_WIDTH : INTEGER := WORD_SIZE);
		PORT(CLK : IN STD_LOGIC;
			  RST : IN STD_LOGIC;
			  EN : IN STD_LOGIC;
			  REG_IN : IN STD_LOGIC_VECTOR(BIT_WIDTH-1 DOWNTO 0);
			  BIT_OUT : OUT STD_LOGIC);
	END COMPONENT;
	COMPONENT COUNTER IS
		GENERIC(BIT_WIDTH : INTEGER := (WORD_SIZE/2+1));
      PORT(CLK : IN STD_LOGIC;
			  RST : IN STD_LOGIC;
           EN : IN STD_LOGIC;
           BITS_OUT : OUT STD_LOGIC_VECTOR(BIT_WIDTH-1 DOWNTO 0));
	END COMPONENT;
	 
	SIGNAL T_FF : STD_LOGIC;
	SIGNAL TOGGLE : STD_LOGIC;
	SIGNAL SHIFT_OUT_SIGNAL : STD_LOGIC;
	SIGNAL SHIFT_IN_SIGNAL : STD_LOGIC;
	SIGNAL DELAY_RESET : STD_LOGIC;
	SIGNAL COUNT_REG : STD_LOGIC_VECTOR(WORD_SIZE/2 DOWNTO 0);
BEGIN
	COUNTER_REG : COUNTER PORT MAP(CLK => CLOCK,
											 RST => NOT T_FF,
											 EN => T_FF,
											 BITS_OUT(WORD_SIZE/2 DOWNTO 0) => COUNT_REG(WORD_SIZE/2 DOWNTO 0));
	MOSI_REG : SHIFT_OUT PORT MAP(CLK => CLOCK, 
											RST => NOT T_FF, 
											EN => NOT SHIFT_OUT_SIGNAL, 
											REG_IN(WORD_SIZE-1 DOWNTO 0) => REG_TX(WORD_SIZE-1 DOWNTO 0), 
											BIT_OUT => MOSI);
	MISO_REG : SHIFT_IN PORT MAP(CLK => CLOCK, 
										  RST => RESET_RX, 
										  EN => SHIFT_IN_SIGNAL, 
										  BIT_IN => MISO, 
										  REG_OUT(WORD_SIZE-1 DOWNTO 0) => REG_RX(WORD_SIZE-1 DOWNTO 0));
	
	SHIFT_IN_SIGNAL <= COUNT_REG(COUNT_REG'HIGH-1);
	SHIFT_OUT_SIGNAL <= (COUNT_REG(2) OR COUNT_REG(1) OR COUNT_REG(0)) AND NOT COUNT_REG(3);
	TOGGLE <= START_TRANSACTION OR DELAY_RESET;
	
	PROCESS(CLOCK)
	BEGIN
		IF CLOCK'EVENT AND CLOCK = '0' THEN
			DELAY_RESET <= COUNT_REG(COUNT_REG'HIGH);
		END IF;
	END PROCESS;

	PROCESS(TOGGLE)
	BEGIN
		IF TOGGLE'EVENT AND TOGGLE = '1' THEN
			T_FF <= NOT T_FF;
		END IF;
	END PROCESS;
	CHIP_SELECT <= NOT T_FF;
END BEHAVIOR;